`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// AUTHOR: ARTHUR J. MILLER
// Create Date: 10/20/2015 05:23:12 PM
// Module Name: Decoder_4to16
// ECE425L LAB #3
// Purpose: 4to16 decoder using 3

// Variables:
//          E : Enable Input
//          S : Selecting Input
//          X = X2X1X0 : 3 bit input  
//          Z : 8 possile outputs, so 8 bit output 

//////////////////////////////////////////////////////////////////////////////////

module Decoder_4to16();
endmodule
