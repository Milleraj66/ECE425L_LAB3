`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// AUTHOR: ARTHUR J. MILLER & Bibek B.
// Module Name: TB_Mux16bit_16to1
// Create Date: 10/20/2015 06:07:50 PM
// ECE425L LAB #3
// Purpose: Develope a Verilog structural model for a 16-bit 16-to-1 MUX
//          Test Bench
//////////////////////////////////////////////////////////////////////////////////

module TB_Mux16bit_16to1();
    // inputs
    reg E;
    reg [3:0] S;
    reg [255:0] X;
    // outputs
    wire [15:0] Z;
    
    // 1. Instatiate Mux module
    //                               Enable,Select(3b),Input0(16b_allIO),Input1,Input2,Input3,Input4,Input5,Input6,Input7, Output
    Mux16bit_16to1       MUX1        (E,S,X,Z);
    
    // 2. Stimulus for test bench
    initial 
        begin
        #5 E=1; S=1;  X[127:112]=128;X[111:96]=64;X[95:80]=32;X[79:64]=16;X[63:48]=8;X[47:32]=4;X[31:16]=2;X[15:0]=1;
        #5 E=1; S=2;  X[127:112]=128;X[111:96]=64;X[95:80]=32;X[79:64]=16;X[63:48]=8;X[47:32]=4;X[31:16]=2;X[15:0]=1;
        #5 E=1; S=3;  X[127:112]=128;X[111:96]=64;X[95:80]=32;X[79:64]=16;X[63:48]=8;X[47:32]=4;X[31:16]=2;X[15:0]=1;
        #5 E=1; S=4;  X[127:112]=128;X[111:96]=64;X[95:80]=32;X[79:64]=16;X[63:48]=8;X[47:32]=4;X[31:16]=2;X[15:0]=1;
        #5 E=1; S=5;  X[127:112]=128;X[111:96]=64;X[95:80]=32;X[79:64]=16;X[63:48]=8;X[47:32]=4;X[31:16]=2;X[15:0]=1;
        #5 E=1; S=6;  X[127:112]=128;X[111:96]=64;X[95:80]=32;X[79:64]=16;X[63:48]=8;X[47:32]=4;X[31:16]=2;X[15:0]=1;
        #5 E=1; S=7;  X[127:112]=128;X[111:96]=64;X[95:80]=32;X[79:64]=16;X[63:48]=8;X[47:32]=4;X[31:16]=2;X[15:0]=1;
        end
endmodule
